`timescale 1ns / 1ps

module model_uart(/*AUTOARG*/
    // Outputs
    TX,
    // Inputs
    RX
    );

    output TX;
    input  RX;

    parameter baud    = 115200;
    parameter bittime = 1000000000/baud;
    parameter name    = "UART0";

    reg [7:0] rxData;
    reg [31:0] rxBuffer; // hold 8 bits
    event     evBit;
    event     evByte;
    event     evTxBit;
    event     evTxByte;
    reg       TX;

    initial
    begin
        TX = 1'b1;
    end

    always @ (negedge RX)
    begin
        rxData[7:0] = 8'h0;
        #(0.5*bittime);

        repeat (8) // 8 bits == 1 byte
        begin
            #bittime ->evBit;
            //rxData[7:0] = {rxData[6:0],RX};
            rxData[7:0] = {RX,rxData[7:1]}; // right shift based on RX bit where RX is the register
        end
        if (rxData[7:0] != 8'h0a && rxData[7:0] != 8'h0d)
        begin
            rxBuffer[31:0] = {rxBuffer[24:0],rxData[7:0]}; // shift by 8
        end
        else
        begin
            if (rxData[7:0] == 8'h0d)
            begin
                $display ("%d %s Received bytes %08x (%s)", $stime, name, rxBuffer, rxBuffer);
            end
        end
        ->evByte;
        // $display ("%d %s Received byte %02x (%s)", $stime, name, rxData, rxData);
    end

    task tskRxData;
    output [7:0] data;
    begin
        @(evByte);
        data = rxData;
    end
    endtask
      
    task tskTxData;
    input [7:0] data;
    reg [9:0]   tmp;
    integer     i;
    begin
        tmp = {1'b1, data[7:0], 1'b0};
        for (i=0;i<10;i=i+1)
        begin
            TX = tmp[i];
            #bittime;
            ->evTxBit;
        end
        ->evTxByte;
    end
    endtask // tskTxData

endmodule // model_uart
