`timescale 1ns / 1ps

module clockCounter(
    input wire in_rst,
    input wire in_norm_clk,
    input wire in_adj_clk,
    input wire in_sel,
    input wire in_adj,
    input wire in_pause,
    output wire [5:0] out_minute,
    output wire [5:0] out_second
    );


endmodule
