`timescale 1ns / 1ps

module snake(
    );

endmodule
